
//frequency lookup table.
//Wavetable has weird register configurations;
//this module is needed to convert piano key frequencies into frequency register contents.
module FrequencyMapper(
	input [4:0] Offset,
	output [23:0] FreqRegValue
);
				
			//25 entries, 24 bit per entry
parameter [0:24][23:0] Freq_ROM = {
	24'b000000011000010011001101,//C4
	24'b000000011001101111101001,//C#4
	24'b000000011011010001101010,//D4
	24'b000000011100111001011100,//D#4
	24'b000000011110100111011011,//E4
	24'b000000100000011011111011,//F4
	24'b000000100010010111011001,//F#4
	24'b000000100100011010001010,//G4
	24'b000000100110100100101010,//G#4
	24'b000000101000110111011111,//A4
	24'b000000101011010010111111,//A#4
	24'b000000101101110111110001,//B4
	24'b000000110000100110011010,//C5
	24'b000000110011011111010010,//C#5
	24'b000000110110100011010100,//D5
	24'b000000111001110010111000,//D#5
	24'b000000111101001110110110,//E5
	24'b000001000000110111110110,//F5
	24'b000001000100101110110010,//F#5
	24'b000001001000110100010100,//G5
	24'b000001001101001001010100,//G#5
	24'b000001010001101110111110,//A5
	24'b000001010110100101111110,//A#5
	24'b000001011011101111100010, //B5
	24'h000000//empty
	};

assign FreqRegValue = Freq_ROM[Offset];

endmodule
