module MIDIFileReader (

);
endmodule
